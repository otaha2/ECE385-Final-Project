module  Frame_control(



							);

							
logic curr_buffer;   //
logic inv_curr_buffer; 






mux2		frame2color(
						.s(inv_curr_buffer),
						.d1(Frame1),
						.d0(Frame0),
						.y()		//output to color mapper
							);

module sprite_table( input logic clk,
							output logic [0:4978][0:23] p1_stand
							
						
							
							);
							

always_comb
begin

p1_stand <=
{
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
32ce2,
2dbc2,
2fc52,
33d22,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
32d22,
30c82,
31cb2,
32d02,
30c72,
2fc42,
2cad2,
23672,
278b2,
30c32,
33d32,
33d42,
32cf2,
30c62,
2fc42,
31ca2,
33d32,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
2fc42,
1f801,
23921,
2cb82,
1d7a1,
18611,
2c693,
697ea,
4a736,
25842,
31cc2,
33d22,
2ab02,
1c711,
18611,
228d1,
32cf2,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
2fc22,
27a11,
2ebf2,
2ec02,
2c922,
3e523,
38613,
2e822,
404d4,
47426,
666b9,
c4c412,
948bd,
455c5,
27941,
269a1,
30833,
394e5,
171e2,
15551,
31cc2,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d32,
32d12,
26971,
10311,
248d1,
248f2,
2f3f3,
ab79b,
89659,
413c4,
b681b,
e4be11,
e9e916,
f7f016,
ecc312,
a277a,
1a231,
101f1,
4f5b8,
a7a910,
4c4b7,
18511,
30c72,
33d22,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d32,
33d32,
30c72,
21871,
3f6d5,
8b93d,
466e6,
455c4,
9c70a,
e49be,
d4a5f,
b39ff,
eaaa10,
ffd514,
fff617,
f4ce13,
aa82c,
7c568,
97679,
9c89c,
baba11,
e3dc15,
b997e,
67616,
1d621,
2aaf2,
33d32,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
2bb22,
27a32,
2bb32,
15551,
52568,
e6e515,
8e7dc,
8c5f9,
eea4f,
ffbf12,
ffde15,
ffed16,
ffbf12,
ffc913,
ffe015,
f2c412,
9c82c,
8875b,
f3bd12,
ffe916,
ffff18,
f5ec16,
cba3f,
6f4c7,
b151 ,
1b6d1,
2bb12,
32d12,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
1b711,
f3e1 ,
248d2,
23572,
645f9,
eee315,
ecbf12,
eba810,
fcbd12,
ffe415,
fff918,
fff016,
ffbf12,
ffb611,
ffc913,
fde816,
eeea16,
ebe716,
fdf417,
fffb18,
ffff18,
e4e115,
786aa,
2f233,
1e1f3,
21333,
27712,
2ebb2,
32cf2,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
33d42,
18631,
3f0  ,
1d3c1,
6e627,
c28ed,
fac312,
ffda15,
ffe516,
ffe816,
fff817,
ffff18,
fff116,
ffbf12,
ffc812,
ffe916,
fffa17,
ffff18,
ffff18,
ffff18,
ffff18,
ffff18,
f3ec16,
c6a0f ,
ac8ad ,
acaa10,
a7a910,
677e9 ,
1e642 ,
2cb72 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
18631 ,
000   ,
1a112 ,
9968a ,
f8a810,
ffaf10,
ffcf14,
ffeb16,
fffc18,
ffff18,
fff217,
ffdf15,
ffd113,
ffe516,
fff918,
ffe916,
fff217,
fffe18,
ffff18,
ffff18,
fff617,
ffe215,
ffd214,
ffdf14,
f5f317,
b7b911,
627c9 ,
1f6b2 ,
2cb92 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
1c741 ,
6190  ,
1b172 ,
9963a ,
f8a310,
fdac11,
e9a722,
e8c325,
fcf41a,
fff617,
f0d020,
deb12c,
dccd31,
dcdc32,
dcd531,
deb52c,
efcf20,
fdef18,
fff317,
fff217,
ffdf15,
ffc712,
ffe216,
f0eb16,
c6c812,
546a7 ,
26752 ,
2ebd2 ,
32d02 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2cb72 ,
1d7b1 ,
212b2 ,
994ea ,
f88c10,
f7a616,
927465,
908e6a,
eee523,
ffd213,
b6924b,
5e5c8f,
536199,
53659a,
536299,
5f5d8e,
b2904e,
f7bd18,
ffc212,
ffc212,
ffbb11,
ffbb11,
ffe516,
b7b711,
46536 ,
2e863 ,
2cb62 ,
32d12 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d32 ,
2db92 ,
28712 ,
5f4c6 ,
8f5224,
93705e,
4a4d9e,
6b6e87,
dabd30,
b5914c,
635a8b,
2136bf,
1932c5,
1932c5,
1932c5,
2237be,
60588d,
947464,
9a7760,
9a7760,
9a7760,
9a7d60,
9a9663,
8a8341,
6a55a ,
356e3 ,
26a02 ,
32cf2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2ebf2 ,
15551 ,
9153e ,
162db8,
1c33c3,
60578e,
b1834d,
4e4d9b,
1831c6,
1c34c5,
283ec2,
3046c4,
364bc8,
364bc9,
364bca,
364bc9,
364bc8,
3046c3,
2c42c1,
2940c1,
1e36c4,
645780,
bf8314,
40314 ,
14521 ,
2bb52 ,
32ce2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32d12 ,
2cb62 ,
13501 ,
9143a ,
162bae,
2134bd,
343fb2,
4348a4,
2639ba,
1831c6,
2d43c0,
7781ad,
a9afba,
c4cad2,
c7cddb,
c8cedf,
c8cedc,
c8ced4,
a8aeba,
9299a8,
7f88a9,
3c4eb4,
263175,
3831b ,
151a1 ,
8230  ,
15591 ,
2cb62 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2dbc2 ,
1b721 ,
a2a0  ,
4a1f  ,
111a5d,
5d4b80,
6354a3,
2336c1,
1831c6,
1831c6,
3448bf,
9499a5,
c7c7aa,
e0e0bf,
f7f7d7,
ffffe3,
ffffe4,
ffffdf,
e9e9c8,
cfcfb0,
a3a498,
414974,
12383d,
19685 ,
1a6b1 ,
1a6b1 ,
1e7f1 ,
2ebf2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2cb72 ,
1f81c ,
e3024 ,
4a14  ,
125   ,
caf   ,
9a6a4b,
b37f7c,
564595,
4f3f98,
494098,
4c4d9c,
7c81a4,
8f95a8,
9aa1b2,
b9c0cb,
c4cada,
c4cade,
c4cadd,
c0c6d3,
aeb2b2,
7c7d72,
2b2c2d,
144e9 ,
2ebf2 ,
30c72 ,
30c72 ,
31ca2 ,
32d22 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
1b701 ,
91c27 ,
10237d,
91146 ,
115   ,
b96   ,
a48451,
e1a262,
ba5f33,
d56327,
c26528,
875946,
4046a1,
2a40c1,
2c42c2,
3147c7,
3349c9,
3349ca,
3349ca,
3248c6,
2a398f,
161929,
775   ,
14501 ,
31cb2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
18641 ,
3613  ,
8103d ,
5923  ,
123   ,
c96   ,
a57445,
f4a05b,
e8843b,
f78d1c,
ee9b2e,
cfa366,
a6a3b4,
545f95,
242661,
7d5c80,
9b6f8a,
9b7e9e,
9ba2ca,
434e85,
7f3d  ,
614c  ,
14531 ,
259b1 ,
32d02 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
1f811 ,
a2c0  ,
6e3   ,
161613,
242420,
2e2922,
a7663b,
ed8948,
f08f45,
fbab35,
ffbe4e,
ffd085,
fcf0c4,
888e91,
36324d,
cc956d,
ffb679,
ffcb95,
fffad4,
6a717e,
7f2e  ,
9219  ,
23922 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2cb52 ,
1d786 ,
152d1b,
474847,
737466,
7d7867,
ad683c,
c85e23,
d06d2d,
f0ac59,
ffbd69,
ffbd7c,
fdebc7,
a0aed9,
5e73cc,
d6cfbf,
ffecb6,
ffefbe,
fff9d6,
8794cb,
293a89,
f291c ,
23922 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
228c1 ,
12421d,
1c3367,
5a607d,
919282,
a6a189,
b57042,
bd5218,
c76023,
ed9854,
ffb86e,
ffcb85,
fef1c2,
dae1db,
c0cbdc,
eff0ce,
fff1b4,
ffe6a3,
ffe5a7,
cebcaa,
7b737a,
203519,
23922 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2fc42 ,
25971 ,
144b24,
c1960 ,
2134a4,
5d6899,
969787,
b3b097,
c8996f,
cc7842,
c55f24,
dd7638,
f29e59,
fdc67e,
ffe7a8,
fef7c1,
fefece,
fffdca,
fff0b3,
ffe199,
ffd786,
edb96d,
a58b43,
3469e ,
29a82 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
28a71 ,
b2c0  ,
e1f62 ,
172fbc,
2239bd,
57639d,
8e908b,
b1b19a,
dcd6b2,
e3bc8e,
c76d37,
c25920,
d97335,
f59e5a,
f9c278,
fce1a1,
fff6c4,
fff6c3,
fff5c1,
fde8ac,
facd7f,
cb8441,
897715,
42b86 ,
32d02 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32d22 ,
28a12 ,
b221  ,
f1b69 ,
1831c6,
1b34c4,
2d42b8,
5763a3,
92948b,
b9b89f,
d6caaa,
e0b893,
ca7441,
c75f25,
d16d31,
d27838,
e7995a,
fdb97c,
fdb97c,
fdb97c,
f1a86a,
d48040,
75431c,
38536 ,
34ba3 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32d12 ,
2aac2 ,
2a703 ,
45308 ,
302a6d,
1831c6,
1831c6,
1831c6,
2e42b8,
5c679c,
8d9093,
babaa3,
dad1b6,
daab84,
d8976b,
d38b5c,
c3612a,
d0672b,
e47e3f,
e47e3f,
e47e3f,
d87d43,
bc7a4c,
4a331e,
10420 ,
2cb62 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32d02 ,
2db62 ,
266c3 ,
42318 ,
9a4513,
734365,
3439b0,
1f33c0,
1831c6,
1a33c5,
233abf,
5c679d,
898e94,
a8aaa9,
d6d2c0,
ece5cb,
e8d2b2,
d08756,
c96929,
cb631b,
cb5f1d,
cb682c,
be7d54,
a09894,
3e3f3d,
10420 ,
2cb62 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d32 ,
2ebe2 ,
1d5d2 ,
4b399 ,
914212,
b74f17,
c45c2a,
a25959,
3c3ca9,
1b32c3,
1a32c4,
1932c5,
2a3fbb,
374ab8,
4b5cb6,
8a8fa1,
b2b3a1,
c9c5ad,
e4d0a9,
eeb660,
f09012,
f07c1d,
eea567,
baa9a8,
4a5ab8,
1a2349,
10420 ,
2cb62 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
29ac2 ,
236b2 ,
4d3b9 ,
873b11,
bd5216,
d75f15,
ef6a12,
e47226,
9c6a5e,
855b71,
62478c,
1f33c0,
1831c6,
1b37cf,
2846d8,
4d64c4,
667ac1,
798ccf,
93a5e0,
cbad7f,
ffa310,
f88320,
c79389,
908bbe,
6a487c,
291d2e,
10420 ,
2cb62 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
20841 ,
191b3 ,
853d11,
be5317,
d46015,
f47811,
fd7810,
fc7e12,
f49819,
f18c1b,
bd6d44,
554f95,
4a44a0,
3e45c0,
2c4ff2,
2d54f8,
3056f8,
3259fa,
375cf9,
977d8a,
f69617,
cf703a,
8a6089,
6a5492,
874028,
3e37c ,
17621 ,
2dbd2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d22 ,
1f7e1 ,
1b123 ,
8e3e12,
d65e15,
f27712,
fd9b10,
ff8910,
ff8010,
ffa110,
ffa710,
f3a019,
dc972c,
d67932,
9c6177,
3d55e8,
2c53fb,
2c53fb,
2c53fb,
2e53f9,
92688a,
dd722c,
704c7f,
78486c,
793d32,
28127 ,
26712 ,
2dbc2 ,
32cf2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
30c62 ,
1f831 ,
374c6 ,
6e32e ,
a74915,
cb5916,
e26a14,
f98711,
ff9010,
ff9110,
ff8e10,
ff8e10,
ff8e10,
ff8e10,
fd9012,
dc8c37,
a58474,
9c837f,
9c837f,
9c7d7f,
9d6b7e,
cc8f7d,
ecab77,
ad6a63,
ab533a,
853b15,
d51   ,
1f811 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2fc42 ,
2a982 ,
35423 ,
7539b ,
c76416,
cc6616,
cc6116,
d45f15,
ea6912,
f88811,
ff9610,
ff7c10,
ff7310,
ff7310,
ff7610,
ff9910,
ffad10,
ffad10,
ffad10,
ffa710,
ff9910,
ff7e12,
ffae5a,
fbd68e,
e88631,
b95512,
6c2fd ,
a41   ,
1f811 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d22 ,
30c62 ,
228c2 ,
253c2 ,
974e9 ,
df77f ,
f29b11,
f39b11,
f38911,
eb7112,
d55f15,
e56c13,
f47610,
ec6cf ,
f56ef ,
fe7310,
ff7510,
ff9510,
ffa710,
ffa810,
ffab10,
ff9b10,
ff8310,
ff7810,
ff9321,
f2a82e,
bb6f1b,
6535c ,
25115 ,
1483  ,
23782 ,
2fc52 ,
32d12 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
30c72 ,
1f812 ,
d370  ,
20162 ,
b652b ,
ff8a10,
ffab10,
ffac10,
ffa210,
f98d10,
e96d12,
de6214,
bd5412,
893da ,
c157c ,
fb7110,
ff7410,
ff8110,
ff8910,
ff8e10,
ffa410,
ffa310,
ff9210,
ff7b10,
ff7e10,
f18111,
b65c15,
5027b ,
2a126 ,
6c2fe ,
3a486 ,
1d7b1 ,
2fc22 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2ebe2 ,
13501 ,
1d172 ,
603d6 ,
ce70d ,
ff9510,
ffaa10,
ff9f10,
ff9910,
fa8d10,
eb6f12,
b14e11,
7432e ,
642ca ,
b551d ,
fa7110,
ff7310,
ff7410,
ff7b10,
ff8b10,
ffa310,
ffac10,
ffa110,
ff7f10,
ff7410,
f77111,
cc5b13,
5d2aa ,
451e7 ,
bf5413,
7739d ,
37436 ,
29892 ,
2ebe2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2dbd2 ,
124b1 ,
54396 ,
e49bf ,
feac10,
ffad10,
ffa710,
ff8310,
ff7410,
f06d12,
c85817,
5a27b ,
2c125 ,
9e4513,
e46613,
fd7210,
ff7310,
ff7410,
ff8710,
ffa710,
ffad10,
ffad10,
ffa210,
ff7f10,
ff7310,
ff7310,
eb6af ,
71337 ,
55265 ,
ed6bf ,
d25d14,
813911,
222b4 ,
23932 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2ebe2 ,
134f1 ,
412d7 ,
ae6f13,
c57d16,
c67e16,
cb8015,
ec8e11,
e77b12,
b35212,
5c28b ,
632bc ,
8a3c11,
b75015,
e46613,
fd7210,
ff7310,
ff7410,
ff7b10,
f98211,
e17813,
d57315,
d56f15,
d46215,
d45e15,
d45e15,
cf5c14,
a54912,
7635d ,
5b296 ,
4a217 ,
2d145 ,
10211 ,
228e1 ,
32d02 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2fc62 ,
1e7d2 ,
2f496 ,
6b4712,
ab6727,
b97026,
ad6918,
cb8214,
af6611,
7436e ,
4d21a ,
853a11,
bd5218,
c45517,
e46613,
fd7210,
ff7410,
ff8010,
ff8110,
f97210,
e06414,
d55e15,
d15c15,
c25417,
bd5218,
c15417,
d05d15,
d56a15,
9851f ,
e71   ,
000   ,
000   ,
4130  ,
165c1 ,
27a32 ,
32d12 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32ce2 ,
2aae2 ,
286f3 ,
4436f ,
bc723d,
db8540,
b26b23,
985c17,
5835b ,
3f1d8 ,
923f12,
b34e17,
c05318,
ca5916,
e36414,
f66f11,
fe7410,
ff8e10,
ff9210,
fe7f10,
fa7a11,
f87911,
ef7312,
d25f16,
c85c17,
cf6216,
e66c13,
f38a11,
af71c ,
11b1  ,
11a3  ,
2018e ,
232419,
111db ,
14521 ,
2aae1 ,
31ca2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2fc42 ,
1a6e1 ,
323d6 ,
805119,
d98545,
f69653,
d28042,
5a3718,
17d3  ,
2e146 ,
a04514,
bd5218,
c85817,
e26414,
db6115,
de6314,
fc7210,
ff7d10,
ff8c10,
ff9c10,
ff9f10,
ff9f10,
fc9510,
f27612,
ee8012,
e98b12,
d86d15,
e98813,
b377b ,
11c1  ,
4c2fd ,
906e3c,
9a9371,
3b3b30,
6150  ,
11450 ,
29a82 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2dbd2 ,
124b1 ,
442912,
be7736,
f1a55c,
ffb56c,
e09f60,
432f1c,
000   ,
1af17 ,
633954,
9b4b3c,
cc5916,
ef6b12,
e96813,
e66713,
fd7110,
ff7410,
ff7e10,
ff9110,
ff9410,
ff9f10,
fa9f10,
e97513,
f07c12,
f38811,
ce6316,
d26f16,
9f5ce ,
f91   ,
663e10,
c18641,
dfb079,
9c714c,
704428,
674923,
356cb ,
27a12 ,
32cf2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2dbd2 ,
124b1 ,
553620,
e4995a,
fec678,
ffd787,
e5c47f,
5f5134,
1612b ,
ff27  ,
2e2e8b,
704269,
af5332,
d0642f,
db6b32,
dc6d35,
de6e34,
ec6e1e,
f46f11,
f46f11,
f46f11,
f48311,
eb8e12,
cb6316,
d96115,
e66917,
b5542c,
a44e33,
753825,
b53   ,
5634d ,
ab6828,
de8a49,
d9864c,
cf7e49,
ba7541,
424615,
1c741 ,
31cb2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2dbd2 ,
124b1 ,
554229,
e6b56f,
ffd383,
ffe29b,
f8e7ac,
cdb176,
695735,
311d16,
803f36,
6c416e,
493c96,
534399,
5c50ad,
6059bc,
655ab6,
a15956,
c4591f,
c55a21,
c55a21,
c55f20,
c1611f,
b95520,
c0571e,
b35732,
5b3f7c,
423996,
342a6b,
d7b   ,
1d104 ,
553311,
965b22,
633c1b,
3b2415,
393113,
2d817 ,
2cb92 ,
32d22 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2dbd2 ,
124b1 ,
553e25,
e6ad6b,
ffdc99,
ffdfa1,
ffcb90,
f6b774,
88633b,
3e20d ,
a04514,
924946,
6b426e,
6c4371,
714c7f,
735289,
735189,
6d477a,
6d477a,
71508a,
72528d,
6e4b80,
6a4272,
6b4270,
906266,
9a715c,
373261,
412f69,
643951,
602b13,
29126 ,
412712,
985c29,
422811,
000   ,
5170  ,
25991 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2dbd2 ,
124b1 ,
432918,
bc7e4f,
f0d39c,
ffd296,
f99d5c,
d0804a,
6b4326,
3a1ba ,
a04514,
bc521a,
ba511b,
bc521b,
c3561b,
c4571b,
b65222,
6a4272,
4341ae,
4a4fc6,
4b52cb,
4547b7,
3f3aa1,
3f399e,
7f6e8e,
a98c68,
553622,
813a12,
c15917,
c86316,
723fc ,
633f18,
975d33,
3e2616,
4110  ,
f3d0  ,
28a51 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2ebf2 ,
14531 ,
12166 ,
423a1d,
b9a066,
f0b874,
d9884e,
604222,
1a158 ,
2e156 ,
a04514,
bd5218,
be5218,
c55617,
df6314,
e26614,
c35919,
ae542b,
a55339,
a7573f,
a75740,
a6553c,
a45137,
a55036,
ca6830,
e47824,
b75817,
ce5d13,
ef7912,
f39a12,
dd90f ,
a46be ,
4a2de ,
1df6  ,
18422 ,
27a11 ,
30c62 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
30ca2 ,
259a1 ,
1d791 ,
27768 ,
566428,
6c5131,
634a23,
3167b ,
10411 ,
2d1b5 ,
a04514,
bd5218,
c55617,
de6314,
f46e11,
f67911,
e58513,
e38613,
e38613,
e38613,
e38613,
e38613,
e38013,
e36d13,
f07c12,
fa9211,
eb8812,
f37c12,
fe8510,
ffa910,
fd9810,
de75e ,
a24ca ,
93429 ,
644c6 ,
1e662 ,
2bb22 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d32 ,
32d02 ,
31cd2 ,
2ebd2 ,
1f6c4 ,
17444 ,
184c3 ,
1f774 ,
16531c,
27253a,
783f48,
8f4d54,
aa594b,
e96e1e,
fe7c10,
fe8a10,
fd9810,
fd9910,
fd9910,
fd9910,
fd9910,
fd9910,
fd9210,
fd7b10,
fe8e10,
fba611,
ee9212,
eb7a12,
f17f12,
fda910,
ff9510,
fd8410,
f88110,
f78010,
b65fb ,
4f385 ,
30792 ,
2bb22 ,
32d12 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32d22 ,
30c62 ,
2dbd2 ,
27a43 ,
1141d ,
d2059 ,
192ca8,
2533b6,
3044d1,
635aba,
d7743e,
fe9618,
ff9b16,
ff7f11,
ff7b10,
ff7a10,
ff7910,
ff7810,
fe7710,
fc7610,
fc7310,
fd8d10,
f49c11,
d06b16,
c35717,
d56e15,
fba410,
ffa710,
ffa610,
ffa710,
ffa810,
f690f ,
d062d ,
46324 ,
19691 ,
31ca2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
269e1 ,
134c10,
102c60,
13279f,
1730c1,
1831c6,
2142e4,
4e62de,
b49589,
eac57f,
fdc866,
fe9c19,
ff9711,
ff8b11,
ff7710,
ff7310,
ee6a12,
d86014,
d65f15,
e97213,
f27e11,
cb5d16,
bd5218,
d06216,
fa8411,
ff8910,
ff9310,
ffa810,
ffad10,
ff9710,
e469e ,
4a285 ,
175e1 ,
30c82 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
1e7f1 ,
4c18  ,
122492,
1831c6,
1933ca,
1d3ad6,
2142e3,
3855de,
7482ba,
9ea7c1,
c1b6a1,
e4b249,
f6be4a,
ffb13a,
ff8a16,
ff7810,
ed6912,
d25c16,
c15417,
b45012,
ad4ed ,
b95115,
bd5218,
ca5816,
e66613,
f66f11,
ff7f10,
ff9410,
ff9a10,
ff8b10,
ea6bf ,
7338a ,
324e5 ,
26952 ,
30c62 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
1e7f1 ,
4c18  ,
122493,
1933ca,
1d3bd7,
254af1,
2d4bde,
384fc6,
4b5ec5,
5567c7,
717bb8,
a49f96,
cac2a9,
e4c585,
f3a431,
fc8116,
fb7111,
e86812,
b14e14,
622bc ,
37185 ,
883b11,
b04c16,
be5317,
c55617,
e36514,
f57011,
f57411,
f57511,
f57311,
ed6a12,
b55113,
5e34c ,
17402 ,
2aaf2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
1e7f1 ,
4c18  ,
122594,
1e3cd9,
2549ef,
2851fc,
5c73d1,
949bb1,
b3baca,
bdc4d1,
97a2ca,
4e5fbc,
5566c3,
8285ac,
c7a36e,
f1842b,
ff7310,
db63e ,
602b9 ,
1cc4  ,
941   ,
35177 ,
813810,
b74f17,
bd5218,
c95817,
d05c16,
d05c16,
d05c16,
d05c16,
ce5b16,
bb5217,
682ed ,
132c1 ,
29a92 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
31ca2 ,
24962 ,
3c5e4 ,
683514,
74455e,
7c558a,
7a5b9a,
6a549f,
917081,
c6976c,
efb87f,
fdc385,
caa793,
6770b2,
6e7dc4,
7885c1,
8581a1,
c48a64,
c06e2e,
844cc ,
32533 ,
c2d0  ,
e62   ,
471f9 ,
8d3d12,
b85017,
bd5218,
bd5218,
be5218,
be5218,
be5218,
be5218,
be5218,
b64f17,
682ed ,
f1b1  ,
19661 ,
29aa1 ,
32d02 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32ce2 ,
2cad2 ,
1e3f1 ,
74347 ,
f87010,
ff7310,
ff7510,
f27112,
cc5f16,
c45a17,
cf5f16,
ee6c12,
f97011,
e68538,
c3b289,
e3d9b2,
b2b2c4,
4d5dbb,
83899b,
616752,
1740a ,
29a92 ,
1d771 ,
221d4 ,
893f11,
ac4a15,
ac4a15,
ac4a15,
ac4b16,
b14c17,
bb5118,
bd5218,
c05318,
c35517,
bd5317,
7736e ,
20132 ,
18101 ,
23682 ,
2ebd2 ,
32d12 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d32 ,
31cd2 ,
289a2 ,
2d4e3 ,
8b4e9 ,
d560d ,
fd7210,
ff7410,
ff8510,
fb9610,
f09512,
ed9412,
e78913,
d76915,
d25e16,
d97620,
e7a435,
f59f42,
d29366,
827f86,
485049,
2e6419,
299e4 ,
30c72 ,
2cb82 ,
28852 ,
323a5 ,
351c7 ,
37187 ,
3d1b8 ,
401c8 ,
662cd ,
ae4c16,
c05618,
d25f15,
eb6c13,
eb6d12,
d673f ,
bc73c ,
b55bb ,
61466 ,
1e601 ,
2ebe2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
31c92 ,
24942 ,
30585 ,
6637b ,
cf5df ,
ff7310,
ff7310,
ff7410,
ff8110,
ff9610,
ffa910,
ffad10,
f7a211,
e38313,
dc6d14,
dd6c14,
e17f14,
f17813,
c66c28,
656240,
2b6317,
23932 ,
31cd2 ,
33d42 ,
33d42 ,
2ec02 ,
1c741 ,
a2d0  ,
1b103 ,
5324b ,
5b27b ,
8139e ,
ca5d13,
dc7414,
ea8312,
fd8e10,
ff8e10,
ff9010,
ff8c10,
f87710,
7c387 ,
17381 ,
2cb62 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2ebf2 ,
15541 ,
42257 ,
b55112,
ed6a11,
ff7310,
ff7410,
ff7d10,
ff8210,
ff8d10,
ffa610,
ffad10,
feac10,
fca410,
fb8e10,
e87313,
c55b16,
c15810,
884fc ,
2c51a ,
29a14 ,
31cc2 ,
33d32 ,
33d42 ,
33d42 ,
32d22 ,
2dbb2 ,
15581 ,
351f6 ,
a54815,
b24d16,
c35615,
e46b13,
ec8612,
ee9412,
f29611,
fb9910,
ff8b10,
ff7810,
f87110,
7c387 ,
17381 ,
2cb62 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2dbd2 ,
124b1 ,
52256 ,
df6410,
fc7111,
ff7310,
ff7910,
ff9710,
ffa510,
ffa610,
ffac10,
ffad10,
ffad10,
ffac10,
ffa710,
ea8b13,
bb5516,
5b2ba ,
284b2 ,
2ca92 ,
31cc2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2fc52 ,
175e1 ,
39217 ,
b04d17,
bd5218,
c05418,
c65717,
c75d17,
c76017,
cd6316,
f07412,
ff7810,
ff7310,
f87010,
7c387 ,
17381 ,
2cb62 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
31ca2 ,
24951 ,
395e3 ,
78428 ,
b55b11,
cf6a14,
cf6e14,
d07f14,
e58912,
fb8d10,
ff8e10,
ff9e10,
ffad10,
ffad10,
ffad10,
cb83e ,
6033b ,
31594 ,
24952 ,
31ca2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
31cd2 ,
269e2 ,
2e614 ,
542bb ,
954013,
bd5218,
bd5218,
bd5218,
cb5817,
e26513,
f76f11,
ff7310,
f87011,
dd6213,
6b2fa ,
16381 ,
2cb62 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d32 ,
269d1 ,
1f452 ,
5e45d ,
975a1b,
b96f27,
bc7127,
d1701d,
e77013,
ea7012,
ea8712,
ee9c11,
fb9f10,
ff9f10,
af6db ,
15151 ,
21891 ,
33d32 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d32 ,
28a42 ,
103d1 ,
5d3ab ,
903f13,
964213,
ab4f16,
ca5f16,
e76e12,
e86e12,
d865f ,
bb55e ,
984411,
4d389 ,
1b5a2 ,
2dbd2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2fc32 ,
26964 ,
203e12,
724b32,
ea9656,
ee9752,
d88239,
ba6a1e,
aa5f16,
a66315,
b56a13,
de7110,
eb74f ,
a254a ,
15201 ,
228f1 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
31ca2 ,
2bb42 ,
25583 ,
21184 ,
311a9 ,
76441b,
a86122,
b96a1d,
b56b1e,
7b4819,
2f1910,
21137 ,
25623 ,
2cb32 ,
32cf2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
28a92 ,
175c13,
173c6f,
75759e,
f8d09b,
fec47e,
efa45c,
bb7437,
593612,
40279 ,
49289 ,
5d2c7 ,
642d6 ,
4e475 ,
247f2 ,
2cb72 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
26a02 ,
15591 ,
f1b12 ,
362f5a,
855d69,
d68745,
d59b54,
816b67,
162060,
5b19  ,
1a6d1 ,
31cb2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32cd2 ,
29ab2 ,
1a6814,
e244d ,
1f3fc7,
6583f1,
c2c9d3,
ebcf98,
dca564,
936b36,
2947a ,
f401  ,
f401  ,
f401  ,
f401  ,
1b6e1 ,
30ca2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32d12 ,
23922 ,
b261e ,
142894,
5b57ba,
b88792,
b99fa3,
777bbd,
2139b8,
c1b59 ,
16531e,
269e4 ,
31cb2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
31ce2 ,
2aaf4 ,
1658f ,
d2349 ,
162ea8,
2244e3,
3257f6,
546fe7,
b3a4a2,
897150,
314612,
2ba03 ,
2dba2 ,
2dba2 ,
2dba2 ,
2dba2 ,
2ec22 ,
32d22 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32d12 ,
23922 ,
c2822 ,
1a33a6,
304fec,
4158e5,
415ce8,
3555ed,
2446e5,
1934bc,
112966,
14491d,
28a66 ,
2dbc2 ,
2fc32 ,
32d02 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d32 ,
2aae2 ,
1656f ,
102e57,
13279c,
1831c2,
1c39d3,
1d3bd8,
2640d4,
4d57b5,
35365e,
1338e ,
2bb32 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32d12 ,
23922 ,
b261f ,
142995,
1d3bd8,
1d3bd8,
1d3bd8,
1d3bd8,
1f3edc,
2244e7,
2040cc,
193b86,
124219,
10440 ,
1a6b1 ,
2dbd2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
28a52 ,
1a6615,
e294c ,
132799,
1831c4,
1831c6,
1831c6,
1831c7,
1932c7,
1a32c2,
152996,
143752,
1d7410,
2aaf2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32d12 ,
23922 ,
92212 ,
a1555 ,
122698,
1832c6,
1d3ad6,
1f3edc,
2943d3,
4d54b3,
6963b3,
72669b,
645746,
615332,
4f6025,
2c859 ,
2cb72 ,
33d22 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
175f2 ,
71134 ,
1429a4,
1831c4,
1832c8,
1934ca,
1a34cb,
1a34cb,
1a34cb,
1a35cc,
2041e0,
1f3fc1,
a1739 ,
1b6db ,
30c62 ,
32d12 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32d12 ,
25982 ,
a2b1  ,
264   ,
9144f ,
1932c4,
2346eb,
274ef9,
3c51d3,
825c58,
bf794c,
e29b6e,
e6bd86,
e6c58b,
aa946c,
2e4026,
20828 ,
2fc42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d22 ,
31cd2 ,
165a6 ,
7e3a  ,
152aa9,
1d33c4,
243dcf,
2b49e5,
2b4de9,
2b4eeb,
2a4eec,
264aed,
2a4ff3,
2d50e9,
2641bb,
193d52,
175f1 ,
2cb82 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d32 ,
2ec12 ,
218a1 ,
b2f0  ,
91249 ,
172fb9,
1b36cb,
1c39d0,
233ac4,
393d9b,
4d4696,
5c57ab,
6470cb,
6675d3,
5265c8,
26429e,
143b3e,
1c735 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2dbd2 ,
20822 ,
134032,
e1d74 ,
2132b0,
594fa7,
7f66a1,
8573b6,
8684c4,
8693d6,
7a92e8,
405ee6,
5165d9,
7f80c7,
8676ba,
3f3656,
c2f0  ,
2aac1 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2cb61 ,
10420 ,
5b2b  ,
d1b6b ,
e1b70 ,
e1b70 ,
e1b70 ,
e1b70 ,
e1b70 ,
102078,
162c8b,
172e90,
172e90,
15297f,
81134 ,
134d4 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
27a31 ,
a280  ,
e2167 ,
162eb9,
2938bb,
816295,
bb7d7b,
bc8482,
bc9c94,
bcb3b1,
a9b3d0,
4d63d4,
6971c1,
b49da5,
c08c90,
5a3f41,
c2f0  ,
2aac1 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
2dbd2 ,
17611 ,
b2e7  ,
d3011 ,
d3012 ,
d3012 ,
d3012 ,
d3012 ,
d3012 ,
d3113 ,
e3316 ,
e3317 ,
e3317 ,
e3214 ,
c2f9  ,
19691 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
269e1 ,
6180  ,
d1c71 ,
1831c6,
1d33c4,
343eb9,
4245b2,
4246b3,
424cb7,
4252bf,
3f55cc,
2f50e8,
395aef,
4d66e8,
5061e2,
262d6a,
c2f0  ,
2aac1 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
32cf2 ,
2db92 ,
29ad2 ,
29ad2 ,
29ad2 ,
29ad2 ,
29ad2 ,
29ad2 ,
29ad2 ,
29ad2 ,
29ad2 ,
29ad2 ,
29ad2 ,
29ad2 ,
29ad2 ,
2dbb2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
269e1 ,
6180  ,
7e38  ,
c1963 ,
c1963 ,
c1963 ,
c1963 ,
c1963 ,
c1963 ,
c1963 ,
d1b65 ,
122577,
15297e,
15297e,
15297e,
a143b ,
c2f0  ,
2aac1 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
29a91 ,
f3c0  ,
a290  ,
a290  ,
a290  ,
a290  ,
a290  ,
a290  ,
a290  ,
a290  ,
a290  ,
a290  ,
a290  ,
a290  ,
a290  ,
a290  ,
134f0 ,
2bb42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
31c92 ,
2aad1 ,
29a91 ,
29a91 ,
29a91 ,
29a91 ,
29a91 ,
29a91 ,
29a91 ,
29a91 ,
29a91 ,
29a91 ,
29a91 ,
29a91 ,
29a91 ,
29a91 ,
2bb22 ,
31cc2 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
33d42 ,
}   
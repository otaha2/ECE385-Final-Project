module player1(input frame_clk 
					
					);
					
					
					